`timescale 1ns/1ps

module cpu_reg (
    input clk,
    input [`DATA_WIDTH-1:0] data_in,
    

);
    
endmodule